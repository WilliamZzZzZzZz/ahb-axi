`ifndef AXI_SEQUENCE_LIB_SV
`define AXI_SEQUENCE_LIB_SV

`include "axi_base_sequence.sv"
`include "axi_master_single_sequence.sv"

`endif